/home/as9397/to_abh/library/Back_End/lef/NangateOpenCellLibrary.lef